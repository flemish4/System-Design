----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    23:23:54 02/06/2018 
-- Design Name: 
-- Module Name:    invRstGen - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity invRstGen is
    Port ( invF : in  STD_LOGIC;
           clk : in  STD_LOGIC;
           invRst : out  STD_LOGIC);
end invRstGen;

architecture Behavioral of invRstGen is
signal invFDelay : std_logic := '0';
begin
	process (clk) begin
		if rising_edge(clk) then
			invFDelay <= invF;
		end if;
	end process;

invRst <= invFDelay and not invF;

end Behavioral;

