`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    03:51:53 02/16/2018 
// Design Name: 
// Module Name:    mux2_8bit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module mux2_8bit(
    input [7:0] A,
    input [7:0] B,
    input SEL,
    output [7:0] X
    );


endmodule
