`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:48:40 01/24/2018 
// Design Name: 
// Module Name:    srl18_8 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module srl18_8(
    input [7:0] D,
    input CE,
    input CLK,
    input [3:0] Addr,
    output [7:0] Q,
    output [7:0] Q15
    );


endmodule
